----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date: 28.09.2022 16:47:14
-- Design Name: Francisco VARELA
-- Module Name: Signal_Generate - Behavioral
-- Project Name:
-- Target Devices:
-- Tool Versions: VERSIO1
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Signal_Generate is
port (clk :in  std_logic;
  --    dataout : out integer range -128 to 127
       --dac_data_o_0 : out std_logic_vector(13 downto 0):=(others => '0')
      -- dac_data_o_0: out std_logic_vector(13 downto 0):=(others => '0')  ;
       dac_sinus_o_0: out std_logic_vector(13 downto 0):=(others => '0') ;
       dac_square_o_0: out std_logic_vector(13 downto 0):=(others => '0')
       );
end Signal_Generate;

architecture Behavioral of Signal_Generate is
signal i : integer range 0 to 2000:=0;
signal signed1 : UNSIGNED(13 downto 0):=(others => '0');
signal signed2 : UNSIGNED(13 downto 0):=(others => '0');
--signal signed1 : UNSIGNED(13 downto 0):=(others => '0');
type memory_type is array (0 to 1999) of integer range 0 to 16384;
--type memory_type is array (0 to 29) of integer range -128 to 127;
--ROM for storing the sine values generated by PYTHON.
--sinus de 2000points
signal sinus: memory_type :=(
8192,8218,8243,8269,8295,8321,8346,8372,8398,8424,8449,8475,8501,8526,8552,8578,8604,8629,8655,8681,8706,8732,8758,8783,8809,8835,8860,8886,8912,8937,8963,8988,9014,9040,9065,9091,9116,9142,9167,9193,9218,9244,9270,9295,9321,9346,9371,9397,9422,9448,9473,9499,9524,9549,9575,9600,9625,9651,9676,9701,9727,9752,9777,9802,9828,9853,9878,9903,9928,9953,9979,10004,10029,10054,10079,10104,10129,10154,10179,10204,10229,10254,10279,10303,10328,10353,10378,10403,10427,10452,10477,10502,10526,10551,10576,10600,10625,10649,10674,10698,10723,
10747,10772,10796,10821,10845,10869,10894,10918,10942,10966,10990,11015,11039,11063,11087,11111,11135,11159,11183,11207,11231,11255,11279,11302,11326,11350,11374,11397,11421,11445,11468,11492,11515,11539,11562,11586,11609,11633,11656,11679,11702,11726,11749,11772,11795,11818,11841,11864,11887,11910,11933,11956,11979,12002,12024,12047,12070,12092,12115,12138,12160,12183,12205,12227,12250,12272,12294,12317,12339,12361,12383,12405,12427,12449,12471,12493,12515,12537,12559,12580,12602,12624,12645,12667,12688,12710,12731,12753,12774,12795,12817,12838,12859,12880,12901,12922,12943,12964,12985,13006,
13027,13047,13068,13089,13109,13130,13150,13171,13191,13212,13232,13252,13272,13293,13313,13333,13353,13373,13393,13413,13432,13452,13472,13491,13511,13531,13550,13569,13589,13608,13627,13647,13666,13685,13704,13723,13742,13761,13780,13798,13817,13836,13854,13873,13892,13910,13928,13947,13965,13983,14001,14019,14038,14056,14073,14091,14109,14127,14145,14162,14180,14197,14215,14232,14250,14267,14284,14301,14318,14335,14352,14369,14386,14403,14420,14436,14453,14470,14486,14503,14519,14535,14551,14568,14584,14600,14616,14632,14648,14663,14679,14695,14710,14726,14741,14757,14772,14787,14803,14818,
14833,14848,14863,14878,14893,14907,14922,14937,14951,14966,14980,14995,15009,15023,15037,15051,15065,15079,15093,15107,15121,15134,15148,15162,15175,15189,15202,15215,15228,15241,15255,15268,15280,15293,15306,15319,15331,15344,15357,15369,15381,15394,15406,15418,15430,15442,15454,15466,15478,15489,15501,15513,15524,15535,15547,15558,15569,15580,15592,15603,15613,15624,15635,15646,15656,15667,15677,15688,15698,15708,15719,15729,15739,15749,15759,15768,15778,15788,15797,15807,15816,15826,15835,15844,15853,15862,15871,15880,15889,15898,15906,15915,15924,15932,15940,15949,15957,15965,15973,15981,
15989,15997,16005,16012,16020,16027,16035,16042,16050,16057,16064,16071,16078,16085,16092,16098,16105,16112,16118,16125,16131,16137,16144,16150,16156,16162,16168,16173,16179,16185,16190,16196,16201,16207,16212,16217,16222,16227,16232,16237,16242,16246,16251,16256,16260,16264,16269,16273,16277,16281,16285,16289,16293,16297,16300,16304,16307,16311,16314,16317,16321,16324,16327,16330,16333,16335,16338,16341,16343,16346,16348,16350,16353,16355,16357,16359,16361,16362,16364,16366,16367,16369,16370,16372,16373,16374,16375,16376,16377,16378,16379,16379,16380,16381,16381,16381,16382,16382,16382,16382,
16382,16382,16382,16381,16381,16381,16380,16379,16379,16378,16377,16376,16375,16374,16373,16372,16370,16369,16367,16366,16364,16362,16361,16359,16357,16355,16353,16350,16348,16346,16343,16341,16338,16335,16333,16330,16327,16324,16321,16317,16314,16311,16307,16304,16300,16297,16293,16289,16285,16281,16277,16273,16269,16264,16260,16256,16251,16246,16242,16237,16232,16227,16222,16217,16212,16207,16201,16196,16190,16185,16179,16173,16168,16162,16156,16150,16144,16137,16131,16125,16118,16112,16105,16098,16092,16085,16078,16071,16064,16057,16050,16042,16035,16027,16020,16012,16005,15997,15989,15981,
15973,15965,15957,15949,15940,15932,15924,15915,15906,15898,15889,15880,15871,15862,15853,15844,15835,15826,15816,15807,15797,15788,15778,15768,15759,15749,15739,15729,15719,15708,15698,15688,15677,15667,15656,15646,15635,15624,15613,15603,15592,15580,15569,15558,15547,15535,15524,15513,15501,15489,15478,15466,15454,15442,15430,15418,15406,15394,15381,15369,15357,15344,15331,15319,15306,15293,15280,15268,15255,15241,15228,15215,15202,15189,15175,15162,15148,15134,15121,15107,15093,15079,15065,15051,15037,15023,15009,14995,14980,14966,14951,14937,14922,14907,14893,14878,14863,14848,14833,14818,
14803,14787,14772,14757,14741,14726,14710,14695,14679,14663,14648,14632,14616,14600,14584,14568,14551,14535,14519,14503,14486,14470,14453,14436,14420,14403,14386,14369,14352,14335,14318,14301,14284,14267,14250,14232,14215,14197,14180,14162,14145,14127,14109,14091,14073,14056,14038,14019,14001,13983,13965,13947,13928,13910,13892,13873,13854,13836,13817,13798,13780,13761,13742,13723,13704,13685,13666,13647,13627,13608,13589,13569,13550,13531,13511,13491,13472,13452,13432,13413,13393,13373,13353,13333,13313,13293,13272,13252,13232,13212,13191,13171,13150,13130,13109,13089,13068,13047,13027,13006,
12985,12964,12943,12922,12901,12880,12859,12838,12817,12795,12774,12753,12731,12710,12688,12667,12645,12624,12602,12580,12559,12537,12515,12493,12471,12449,12427,12405,12383,12361,12339,12317,12294,12272,12250,12227,12205,12183,12160,12138,12115,12092,12070,12047,12024,12002,11979,11956,11933,11910,11887,11864,11841,11818,11795,11772,11749,11726,11702,11679,11656,11633,11609,11586,11562,11539,11515,11492,11468,11445,11421,11397,11374,11350,11326,11302,11279,11255,11231,11207,11183,11159,11135,11111,11087,11063,11039,11015,10990,10966,10942,10918,10894,10869,10845,10821,10796,10772,10747,10723,
10698,10674,10649,10625,10600,10576,10551,10526,10502,10477,10452,10427,10403,10378,10353,10328,10303,10279,10254,10229,10204,10179,10154,10129,10104,10079,10054,10029,10004,9979,9953,9928,9903,9878,9853,9828,9802,9777,9752,9727,9701,9676,9651,9625,9600,9575,9549,9524,9499,9473,9448,9422,9397,9371,9346,9321,9295,9270,9244,9218,9193,9167,9142,9116,9091,9065,9040,9014,8988,8963,8937,8912,8886,8860,8835,8809,8783,8758,8732,8706,8681,8655,8629,8604,8578,8552,8526,8501,8475,8449,8424,8398,8372,8346,8321,8295,8269,8243,8218,8192,
8166,8141,8115,8089,8063,8038,8012,7986,7960,7935,7909,7883,7858,7832,7806,7780,7755,7729,7703,7678,7652,7626,7601,7575,7549,7524,7498,7472,7447,7421,7396,7370,7344,7319,7293,7268,7242,7217,7191,7166,7140,7114,7089,7063,7038,7013,6987,6962,6936,6911,6885,6860,6835,6809,6784,6759,6733,6708,6683,6657,6632,6607,6582,6556,6531,6506,6481,6456,6431,6405,6380,6355,6330,6305,6280,6255,6230,6205,6180,6155,6130,6105,6081,6056,6031,6006,5981,5957,5932,5907,5882,5858,5833,5808,5784,5759,5735,5710,5686,5661,
5637,5612,5588,5563,5539,5515,5490,5466,5442,5418,5394,5369,5345,5321,5297,5273,5249,5225,5201,5177,5153,5129,5105,5082,5058,5034,5010,4987,4963,4939,4916,4892,4869,4845,4822,4798,4775,4751,4728,4705,4682,4658,4635,4612,4589,4566,4543,4520,4497,4474,4451,4428,4405,4382,4360,4337,4314,4292,4269,4246,4224,4201,4179,4157,4134,4112,4090,4067,4045,4023,4001,3979,3957,3935,3913,3891,3869,3847,3825,3804,3782,3760,3739,3717,3696,3674,3653,3631,3610,3589,3567,3546,3525,3504,3483,3462,3441,3420,3399,3378,
3357,3337,3316,3295,3275,3254,3234,3213,3193,3172,3152,3132,3112,3091,3071,3051,3031,3011,2991,2971,2952,2932,2912,2893,2873,2853,2834,2815,2795,2776,2757,2737,2718,2699,2680,2661,2642,2623,2604,2586,2567,2548,2530,2511,2492,2474,2456,2437,2419,2401,2383,2365,2346,2328,2311,2293,2275,2257,2239,2222,2204,2187,2169,2152,2134,2117,2100,2083,2066,2049,2032,2015,1998,1981,1964,1948,1931,1914,1898,1881,1865,1849,1833,1816,1800,1784,1768,1752,1736,1721,1705,1689,1674,1658,1643,1627,1612,1597,1581,1566,
1551,1536,1521,1506,1491,1477,1462,1447,1433,1418,1404,1389,1375,1361,1347,1333,1319,1305,1291,1277,1263,1250,1236,1222,1209,1195,1182,1169,1156,1143,1129,1116,1104,1091,1078,1065,1053,1040,1027,1015,1003,990,978,966,954,942,930,918,906,895,883,871,860,849,837,826,815,804,792,781,771,760,749,738,728,717,707,696,686,676,665,655,645,635,625,616,606,596,587,577,568,558,549,540,531,522,513,504,495,486,478,469,460,452,444,435,427,419,411,403,
395,387,379,372,364,357,349,342,334,327,320,313,306,299,292,286,279,272,266,259,253,247,240,234,228,222,216,211,205,199,194,188,183,177,172,167,162,157,152,147,142,138,133,128,124,120,115,111,107,103,99,95,91,87,84,80,77,73,70,67,63,60,57,54,51,49,46,43,41,38,36,34,31,29,27,25,23,22,20,18,17,15,14,12,11,10,9,8,7,6,5,5,4,3,3,3,0,0,0,0,
0,0,0,3,3,3,4,5,5,6,7,8,9,10,11,12,14,15,17,18,20,22,23,25,27,29,31,34,36,38,41,43,46,49,51,54,57,60,63,67,70,73,77,80,84,87,91,95,99,103,107,111,115,120,124,128,133,138,142,147,152,157,162,167,172,177,183,188,194,199,205,211,216,222,228,234,240,247,253,259,266,272,279,286,292,299,306,313,320,327,334,342,349,357,364,372,379,387,395,403,
411,419,427,435,444,452,460,469,478,486,495,504,513,522,531,540,549,558,568,577,587,596,606,616,625,635,645,655,665,676,686,696,707,717,728,738,749,760,771,781,792,804,815,826,837,849,860,871,883,895,906,918,930,942,954,966,978,990,1003,1015,1027,1040,1053,1065,1078,1091,1104,1116,1129,1143,1156,1169,1182,1195,1209,1222,1236,1250,1263,1277,1291,1305,1319,1333,1347,1361,1375,1389,1404,1418,1433,1447,1462,1477,1491,1506,1521,1536,1551,1566,
1581,1597,1612,1627,1643,1658,1674,1689,1705,1721,1736,1752,1768,1784,1800,1816,1833,1849,1865,1881,1898,1914,1931,1948,1964,1981,1998,2015,2032,2049,2066,2083,2100,2117,2134,2152,2169,2187,2204,2222,2239,2257,2275,2293,2311,2328,2346,2365,2383,2401,2419,2437,2456,2474,2492,2511,2530,2548,2567,2586,2604,2623,2642,2661,2680,2699,2718,2737,2757,2776,2795,2815,2834,2853,2873,2893,2912,2932,2952,2971,2991,3011,3031,3051,3071,3091,3112,3132,3152,3172,3193,3213,3234,3254,3275,3295,3316,3337,3357,3378,
3399,3420,3441,3462,3483,3504,3525,3546,3567,3589,3610,3631,3653,3674,3696,3717,3739,3760,3782,3804,3825,3847,3869,3891,3913,3935,3957,3979,4001,4023,4045,4067,4090,4112,4134,4157,4179,4201,4224,4246,4269,4292,4314,4337,4360,4382,4405,4428,4451,4474,4497,4520,4543,4566,4589,4612,4635,4658,4682,4705,4728,4751,4775,4798,4822,4845,4869,4892,4916,4939,4963,4987,5010,5034,5058,5082,5105,5129,5153,5177,5201,5225,5249,5273,5297,5321,5345,5369,5394,5418,5442,5466,5490,5515,5539,5563,5588,5612,5637,5661,
5686,5710,5735,5759,5784,5808,5833,5858,5882,5907,5932,5957,5981,6006,6031,6056,6081,6105,6130,6155,6180,6205,6230,6255,6280,6305,6330,6355,6380,6405,6431,6456,6481,6506,6531,6556,6582,6607,6632,6657,6683,6708,6733,6759,6784,6809,6835,6860,6885,6911,6936,6962,6987,7013,7038,7063,7089,7114,7140,7166,7191,7217,7242,7268,7293,7319,7344,7370,7396,7421,7447,7472,7498,7524,7549,7575,7601,7626,7652,7678,7703,7729,7755,7780,7806,7832,7858,7883,7909,7935,7960,7986,8012,8038,8063,8089,8115,8141,8166
);
--60pontos
--signal square0 :memory_type:=(16382 , 16382 , 16382 , 16382 ,
--16382 , 16382 , 16382 , 16382 , 16382 , 16382 ,
--16382 , 16382 , 16382 , 16382 , 16382 , 16382 ,
--16382 , 16382 , 16382 , 16382 , 16382 , 16382 ,
--16382 , 16382 , 16382 , 16382 , 16382 , 16382 ,
-- 16382 , 16382 , 2 , 2 , 2 , 2 , 2 , 2 , 2,
-- 2 , 2 , 2 , 2 , 2 , 2 , 2 , 2 , 2 , 2 , 2 , 2 , 2 ,
-- 2 , 2 , 2 , 2 , 2 , 2 , 2 , 2 , 2 , 2  );
-- --60pontos
-- signal square10 :memory_type:=(16382 , 16382 , 16382 , 16382 ,
--16382 , 16382 , 16382 , 16382 , 16382 , 16382 ,
--16382 , 16382 , 16382 , 16382 , 16382 , 16382 ,
--16382 , 16382 , 16382 , 16382 , 16382 , 16382 ,
--16382 , 16382 , 16382 , 16382 , 16382 , 8192,
--8192 ,8192 , 2 , 2 , 2 , 2 , 2 , 2 , 2,
-- 2 , 2 , 2 , 2 , 2 , 2 , 2 , 2 , 2 , 2 , 2 , 2 , 2 ,
-- 2 , 2 , 2 , 2 , 2 , 2 , 2 , 8192 ,8192 ,8192  );
 --2000pontos
 signal square0_2000 :memory_type:=(16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0
);
signal square10_2000 :memory_type:=(16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192
);

signal square15_2000 :memory_type:=(
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192
);

signal square50_2000 :memory_type:=(
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,
16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,16382,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,
0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,
8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192,8192
);
--signal sine : memory_type :=(9540, 12296, 14204, 15688, 16324, 16324, 15688, 14204, 12296, 9540); --, -3392, -6572, -9540, -12296, -14204, -15688, -16324, -16324, -15688, -14204, -12296, -9540, -6572, -3392
--ORIGINal
--signal sine : memory_type :=(0, 3392, 6572, 9540, 12296, 14204, 15688, 16324, 16324, 15688, 14204, 12296, 9540,
--6572, 3392, -3392, -6572, -9540, -12296, -14204, -15688, -16324, -16324, -15688, -14204, -12296, -9540, -6572, -3392
--original
--signal sine : memory_type :=(0,16,31,45,58,67,74,77,77,74,67,58,45,31,16,0,
---16,-31,-45,-58,-67,-74,-77,-77,-74,-67,-58,-45,-31,-16);
begin

process(clk)
begin
  --to check the rising edge of the clock signal
if(rising_edge(clk)) then
--dataout <= sine(i);
--signed1 <= TO_UNSIGNED(sine(i),14);
signed1 <= TO_UNSIGNED(sinus(i),14);
signed2 <= TO_UNSIGNED(square15_2000(i),14);
dac_sinus_o_0<= STD_LOGIC_VECTOR(signed1);
dac_square_o_0<= STD_LOGIC_VECTOR(signed2);
i <= i+ 1;
if(i = 1999) then
i <= 0;
end if;
end if;
end process;

end Behavioral;